// Testbench for cpu module