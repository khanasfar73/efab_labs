module regfile(
        rd_addr, wr_addr, rd_data, wr_data
    );

endmodule
