// Top module for the CPU core

module cpu();
    // TODO
endmodule
